`timescale 1ns / 1ps

module ntt_const_lut(
    input forward,
    input [7:0] idx,
    output reg [63:0] val
);

always @(forward, idx) begin
    case ({~forward, idx}) // TODO improve
        9'h000: val <= 64'h7b14d0c689871ae6;
        9'h001: val <= 64'h23aadfb5edf35d70;
        9'h002: val <= 64'h111abd573830ef07;
        9'h003: val <= 64'hf821f1b771202bcb;
        9'h004: val <= 64'had2d23357a5ddaa3;
        9'h005: val <= 64'h1e365b58f203fd54;
        9'h006: val <= 64'h91103a3e12ecae09;
        9'h007: val <= 64'h5de6e61530f1d512;
        9'h008: val <= 64'haa0bbfca2de3d915;
        9'h009: val <= 64'hfd657fa55a4c81b6;
        9'h00a: val <= 64'h6804c8e77418e117;
        9'h00b: val <= 64'h6172322940eba85d;
        9'h00c: val <= 64'he7dc1787cf78533b;
        9'h00d: val <= 64'h57a6bc1220e4198e;
        9'h00e: val <= 64'hae19ca2e4f30ebce;
        9'h00f: val <= 64'hcb535a60ede2b6bd;
        9'h010: val <= 64'hd0096bbd202dc3e4;
        9'h011: val <= 64'h0258076723f5dbc4;
        9'h012: val <= 64'h9ef9e03fa16485b4;
        9'h013: val <= 64'h891ba983e4c88a87;
        9'h014: val <= 64'hc396831a77d55dda;
        9'h015: val <= 64'hc651d94cf106169c;
        9'h016: val <= 64'h2a56599274c87bea;
        9'h017: val <= 64'h7d9344fcbdbe2d3c;
        9'h018: val <= 64'hb495f7375776e5b6;
        9'h019: val <= 64'h552165817f4b4912;
        9'h01a: val <= 64'h629cff70e6ab2f95;
        9'h01b: val <= 64'haed76417a41a4c00;
        9'h01c: val <= 64'h4d68443ac0f5960d;
        9'h01d: val <= 64'h8ec5a11fb226cf46;
        9'h01e: val <= 64'h770b56e9744edbc0;
        9'h01f: val <= 64'h5b7d3dc41a830f86;
        9'h020: val <= 64'h9a0624b721b31403;
        9'h021: val <= 64'h533a47a03f370097;
        9'h022: val <= 64'h4500b4ebc56124cf;
        9'h023: val <= 64'ha3b59cbffcaf29ee;
        9'h024: val <= 64'h3e6a18ab3332eb39;
        9'h025: val <= 64'h5bf29bd34ca5c72e;
        9'h026: val <= 64'he2354362b5054065;
        9'h027: val <= 64'hb0cbed29fd63ec75;
        9'h028: val <= 64'h28687d52c24d8a9b;
        9'h029: val <= 64'h932296f3c07a1ffd;
        9'h02a: val <= 64'h44ead90859d57b34;
        9'h02b: val <= 64'hf8a416df3a1ce3e9;
        9'h02c: val <= 64'hf2b36b56d2a614e3;
        9'h02d: val <= 64'hc7b35de8fea7219c;
        9'h02e: val <= 64'hd5f715a2bfedaeca;
        9'h02f: val <= 64'h43192ea1785957ab;
        9'h030: val <= 64'h8ce09165945ad1ba;
        9'h031: val <= 64'h9cfca3e3f424ab9b;
        9'h032: val <= 64'h62648df161c96353;
        9'h033: val <= 64'hf1cbe173c176f96d;
        9'h034: val <= 64'h3fc5d9f5eb6d8e9b;
        9'h035: val <= 64'h1286ad4a2534e675;
        9'h036: val <= 64'h35204479dc9da5fd;
        9'h037: val <= 64'hd4b3c7bfb42b8bb9;
        9'h038: val <= 64'hbd49348cd79bbfab;
        9'h039: val <= 64'h2bac8ea2abdb41a4;
        9'h03a: val <= 64'he6e09ac4ab930600;
        9'h03b: val <= 64'h556dea00a29198f8;
        9'h03c: val <= 64'hf3819f473ba4753b;
        9'h03d: val <= 64'hd646737b6bb09af9;
        9'h03e: val <= 64'h13edf74417ea2fd1;
        9'h03f: val <= 64'h3dd4da460cc97d4a;
        9'h040: val <= 64'h25edb38ab4bd5053;
        9'h041: val <= 64'hd6e7d01a34f0a811;
        9'h042: val <= 64'hd7b7a85190f81a3b;
        9'h043: val <= 64'h75e05007850f0083;
        9'h044: val <= 64'h7c87cea914f50b00;
        9'h045: val <= 64'ha122bc70ba22d39f;
        9'h046: val <= 64'h93cb97c2ef88ee0d;
        9'h047: val <= 64'h52d0ee647eafba09;
        9'h048: val <= 64'h90fb7c5d0a31ea27;
        9'h049: val <= 64'hb97b4d1b6def702d;
        9'h04a: val <= 64'h0bc9612c124e8e9a;
        9'h04b: val <= 64'h29dc4ddac558c74c;
        9'h04c: val <= 64'h5381d29a568de781;
        9'h04d: val <= 64'h523ecb16d8fa59fa;
        9'h04e: val <= 64'h6b78f0610a714386;
        9'h04f: val <= 64'h01839215423cecec;
        9'h050: val <= 64'hd045b507156a83dd;
        9'h051: val <= 64'h747fa042d0127ec3;
        9'h052: val <= 64'h81a8a6090d936c84;
        9'h053: val <= 64'hbc977d3d8a12df28;
        9'h054: val <= 64'h13028e6629130438;
        9'h055: val <= 64'h29a912834df1e37e;
        9'h056: val <= 64'h960978f89984a7fb;
        9'h057: val <= 64'hc3b3bda8b90ae584;
        9'h058: val <= 64'hf4b71741e67dced2;
        9'h059: val <= 64'hb3f6b5d3f637f7e6;
        9'h05a: val <= 64'h86d97dd7038637f7;
        9'h05b: val <= 64'h07590e9403f2ff42;
        9'h05c: val <= 64'hf38b1dd44a359469;
        9'h05d: val <= 64'h1f7241c1961b6c25;
        9'h05e: val <= 64'h0820e364b164b241;
        9'h05f: val <= 64'h495d36ba9ab2221a;
        9'h060: val <= 64'h58610d63888e6bbb;
        9'h061: val <= 64'h020716534aa1ba32;
        9'h062: val <= 64'had851115167dcd9e;
        9'h063: val <= 64'heef4c8f716f0de87;
        9'h064: val <= 64'h841db197137d9e93;
        9'h065: val <= 64'h3e6fbad13f00422e;
        9'h066: val <= 64'hc1668bda4bccf8af;
        9'h067: val <= 64'h3db0a40daea26322;
        9'h068: val <= 64'h499ed16d6696670a;
        9'h069: val <= 64'h9f5ed952badd057f;
        9'h06a: val <= 64'h73c50fd40f3a4264;
        9'h06b: val <= 64'h2b25e6840a99de53;
        9'h06c: val <= 64'h7bb618d11368aa4f;
        9'h06d: val <= 64'h2a1057cbcccee8a3;
        9'h06e: val <= 64'h741e6c2cb6da9491;
        9'h06f: val <= 64'h6e5704bab42410ec;
        9'h070: val <= 64'h2ccb2b30a74f74ba;
        9'h071: val <= 64'ha4a0dfe61f56f176;
        9'h072: val <= 64'h555f30304de95af0;
        9'h073: val <= 64'h43ff75349014b293;
        9'h074: val <= 64'h149c337155c30125;
        9'h075: val <= 64'h455d9d591d2db1c3;
        9'h076: val <= 64'h963793afcf9fe50a;
        9'h077: val <= 64'hac95d15f1765532b;
        9'h078: val <= 64'he9c1f2424d1e196c;
        9'h079: val <= 64'h0fa3f9ca176c4c13;
        9'h07a: val <= 64'hebc3fd84163a5cfc;
        9'h07b: val <= 64'hdf3ec3908447746c;
        9'h07c: val <= 64'h0d4fef6a64b3fe7b;
        9'h07d: val <= 64'h3e145968b25ab326;
        9'h07e: val <= 64'h824d345592851bf8;
        9'h07f: val <= 64'h00a93c121c10b0af;
        9'h080: val <= 64'h59a8473ba280634b;
        9'h081: val <= 64'hb9067dc2d63720b6;
        9'h082: val <= 64'hf683298843ed4555;
        9'h083: val <= 64'h46ffc5af9e9a6032;
        9'h084: val <= 64'h8d601c135df9e29d;
        9'h085: val <= 64'h41d7046590d01d53;
        9'h086: val <= 64'he94aa030f45c27ec;
        9'h087: val <= 64'hab4f216aca169db1;
        9'h088: val <= 64'hcdcc7796ee798973;
        9'h089: val <= 64'h794976ba2654bc62;
        9'h08a: val <= 64'hd7ad3433540e63a5;
        9'h08b: val <= 64'h1323c7e126c9839a;
        9'h08c: val <= 64'h3bca582585db15b7;
        9'h08d: val <= 64'h857b375b4f60af2c;
        9'h08e: val <= 64'h6d8b12985da00e5d;
        9'h08f: val <= 64'h6d506698e206e63e;
        9'h090: val <= 64'h577967387b179fad;
        9'h091: val <= 64'h0b639aeaaa499ba7;
        9'h092: val <= 64'h583e76a5c837779c;
        9'h093: val <= 64'h6bf62b30794ff2a7;
        9'h094: val <= 64'h3ce2456885f823ae;
        9'h095: val <= 64'h6dd489ae9fdc4e94;
        9'h096: val <= 64'hf9c4302418846559;
        9'h097: val <= 64'h240f6001ef69a6ca;
        9'h098: val <= 64'hc40658f32c0a2f70;
        9'h099: val <= 64'ha0db14725879d89a;
        9'h09a: val <= 64'h4296db5f3aa2baab;
        9'h09b: val <= 64'h29fa75db424a74a5;
        9'h09c: val <= 64'h2aadc5fc1fd685d6;
        9'h09d: val <= 64'he876962d7a571e64;
        9'h09e: val <= 64'hfc4de89fda39ae89;
        9'h09f: val <= 64'h82318159db77680d;
        9'h0a0: val <= 64'he23a0cbae4129738;
        9'h0a1: val <= 64'h947df33e69abfa91;
        9'h0a2: val <= 64'hfb067124e287466f;
        9'h0a3: val <= 64'hba8ce07e9f221f57;
        9'h0a4: val <= 64'ha3e50a7b5ffddc5f;
        9'h0a5: val <= 64'hca60de75bddb51f1;
        9'h0a6: val <= 64'hfb01c7db0fe39956;
        9'h0a7: val <= 64'h8e9a9d420d594b7f;
        9'h0a8: val <= 64'h2c53a3914388ed62;
        9'h0a9: val <= 64'hbd780b839ee787bf;
        9'h0aa: val <= 64'h859f2c14a7ef75ec;
        9'h0ab: val <= 64'hb542fd5a463b9030;
        9'h0ac: val <= 64'h3e7e644cf61cf72e;
        9'h0ad: val <= 64'h68d3f1127653d1c0;
        9'h0ae: val <= 64'h5aefcb7c711a0727;
        9'h0af: val <= 64'h4a2816b2ea29ebad;
        9'h0b0: val <= 64'hcedcf34e539af2c0;
        9'h0b1: val <= 64'h80a085795ddc7d09;
        9'h0b2: val <= 64'he95c7abc0589ef7f;
        9'h0b3: val <= 64'h5c2f6ed927f75242;
        9'h0b4: val <= 64'h7971c9eddabe1e75;
        9'h0b5: val <= 64'h4898689f6fc23f00;
        9'h0b6: val <= 64'h3bbdbe33c55dd1bf;
        9'h0b7: val <= 64'h745a97b0851c0641;
        9'h0b8: val <= 64'hfd31be61c01063b9;
        9'h0b9: val <= 64'h3f01e5b34fae0aa7;
        9'h0ba: val <= 64'h7e189ce17128ea7f;
        9'h0bb: val <= 64'h781fc1e2cb388266;
        9'h0bc: val <= 64'h71ac19188eb4a196;
        9'h0bd: val <= 64'h439aced2e3b95ca6;
        9'h0be: val <= 64'h5b76829a7d312b48;
        9'h0bf: val <= 64'h966daa7acdf136e8;
        9'h0c0: val <= 64'h0356aa26a444769f;
        9'h0c1: val <= 64'h75230cecaf71b841;
        9'h0c2: val <= 64'hd72e468d985d555c;
        9'h0c3: val <= 64'h461fa87b1166a135;
        9'h0c4: val <= 64'ha2f46adfb3e8142f;
        9'h0c5: val <= 64'h1bf20b7597280162;
        9'h0c6: val <= 64'hbf6a7c11d2de0a24;
        9'h0c7: val <= 64'h1d353167326aba7c;
        9'h0c8: val <= 64'hd0f012076961cf97;
        9'h0c9: val <= 64'h1c8f7a522126036d;
        9'h0ca: val <= 64'hcf8889e072edeeb3;
        9'h0cb: val <= 64'h55dae99cca9f43d2;
        9'h0cc: val <= 64'hd15063bb94572a61;
        9'h0cd: val <= 64'hce4131c5343f1195;
        9'h0ce: val <= 64'h34679e4f84b49624;
        9'h0cf: val <= 64'hc0409a0bc48c1336;
        9'h0d0: val <= 64'hda592af687a0bf83;
        9'h0d1: val <= 64'he94a2e84ebac033d;
        9'h0d2: val <= 64'ha0fd4342d733010b;
        9'h0d3: val <= 64'h093ee1cee28b5fb3;
        9'h0d4: val <= 64'h8b22c29915c2a850;
        9'h0d5: val <= 64'h9f7617ab77c9d9e6;
        9'h0d6: val <= 64'h6d779b0f82f63cd5;
        9'h0d7: val <= 64'he58d75de55cd6ba5;
        9'h0d8: val <= 64'h363cf96d96b48aae;
        9'h0d9: val <= 64'he9cc7798d1a1d61d;
        9'h0da: val <= 64'h0be985c732f3a244;
        9'h0db: val <= 64'h8e07006b8aaa770f;
        9'h0dc: val <= 64'hb4d7601889758cd3;
        9'h0dd: val <= 64'h86f6dc87dc59ebdc;
        9'h0de: val <= 64'h94705fb38d84dfec;
        9'h0df: val <= 64'h9f7068937866b200;
        9'h0e0: val <= 64'h3200b7cec5fe17f3;
        9'h0e1: val <= 64'ha9239fde2cd60394;
        9'h0e2: val <= 64'h077063a6dac6fc5d;
        9'h0e3: val <= 64'h5c1a64c06b7dd046;
        9'h0e4: val <= 64'h289a3925f94c8124;
        9'h0e5: val <= 64'ha6c6de29adaf173e;
        9'h0e6: val <= 64'h13f8105c8a951ed3;
        9'h0e7: val <= 64'h812ec865d84ea283;
        9'h0e8: val <= 64'h8e17933de1837acb;
        9'h0e9: val <= 64'h70411dccc13d8b61;
        9'h0ea: val <= 64'h4289f6df6059e2f7;
        9'h0eb: val <= 64'h3fa72e9cb12ca689;
        9'h0ec: val <= 64'h64b8908e5bd418f7;
        9'h0ed: val <= 64'h1cb446215d95bd16;
        9'h0ee: val <= 64'h1ca69e37838cdded;
        9'h0ef: val <= 64'h4f0831687b9a69a0;
        9'h0f0: val <= 64'h586702a02334ebf8;
        9'h0f1: val <= 64'h6c904e3d6aeec005;
        9'h0f2: val <= 64'h22256ef5c744e616;
        9'h0f3: val <= 64'hf97e2b576eca967c;
        9'h0f4: val <= 64'hfa4c2a463c91553b;
        9'h0f5: val <= 64'hbb1ccfc281bf5233;
        9'h0f6: val <= 64'h2970df9aeaf9d2fc;
        9'h0f7: val <= 64'h87e645caf2b023a5;
        9'h0f8: val <= 64'ha0f1c104e7d2a04a;
        9'h0f9: val <= 64'h833a08a8290e0029;
        9'h0fa: val <= 64'h9f8ae77d6e7aa38c;
        9'h0fb: val <= 64'hf54b1db3d9c1a7cf;
        9'h0fc: val <= 64'he31abb31fc784aab;
        9'h0fd: val <= 64'h674eb812226a87a4;
        9'h0fe: val <= 64'h1f9b744f63af4b31;
        // backward
        9'h100: val <= 64'he03a2942eba63cd0;
        9'h101: val <= 64'h9886e5802ceb005d;
        9'h102: val <= 64'h1cbae26052dd3d56;
        9'h103: val <= 64'h0a8a7fde7593e032;
        9'h104: val <= 64'h604ab614e0dae475;
        9'h105: val <= 64'h7c9b94ea264787d8;
        9'h106: val <= 64'h5ee3dc8d6782e7b7;
        9'h107: val <= 64'h77ef57c75ca5645c;
        9'h108: val <= 64'hd664bdf7645bb505;
        9'h109: val <= 64'h44b8cdcfcd9635ce;
        9'h10a: val <= 64'h0589734c12c432c6;
        9'h10b: val <= 64'h0657723ae08af185;
        9'h10c: val <= 64'hddb02e9c8810a1eb;
        9'h10d: val <= 64'h93454f54e466c7fc;
        9'h10e: val <= 64'ha76e9af22c209c09;
        9'h10f: val <= 64'hb0cd6c29d3bb1e61;
        9'h110: val <= 64'he32eff5acbc8aa14;
        9'h111: val <= 64'he3215770f1bfcaeb;
        9'h112: val <= 64'h9b1d0d03f3816f0a;
        9'h113: val <= 64'hc02e6ef59e28e178;
        9'h114: val <= 64'hbd4ba6b2eefba50a;
        9'h115: val <= 64'h8f947fc58e17fca0;
        9'h116: val <= 64'h71be0a546dd20d36;
        9'h117: val <= 64'h7ea6d52c7706e57e;
        9'h118: val <= 64'hebdd8d35c4c0692e;
        9'h119: val <= 64'h590ebf68a1a670c3;
        9'h11a: val <= 64'hd73b646c560906dd;
        9'h11b: val <= 64'ha3bb38d1e3d7b7bb;
        9'h11c: val <= 64'hf86539eb748e8ba4;
        9'h11d: val <= 64'h56b1fdb4227f846d;
        9'h11e: val <= 64'hcdd4e5c38957700e;
        9'h11f: val <= 64'h606534fed6eed601;
        9'h120: val <= 64'h6b653ddec1d0a815;
        9'h121: val <= 64'h78dec10a72fb9c25;
        9'h122: val <= 64'h4afe3d79c5dffb2e;
        9'h123: val <= 64'h71ce9d26c4ab10f2;
        9'h124: val <= 64'hf3ec17cb1c61e5bd;
        9'h125: val <= 64'h160925f97db3b1e4;
        9'h126: val <= 64'hc998a424b8a0fd53;
        9'h127: val <= 64'h1a4827b3f9881c5c;
        9'h128: val <= 64'h925e0282cc5f4b2c;
        9'h129: val <= 64'h605f85e6d78bae1b;
        9'h12a: val <= 64'h74b2daf93992dfb1;
        9'h12b: val <= 64'hf696bbc36cca284e;
        9'h12c: val <= 64'h5ed85a4f782286f6;
        9'h12d: val <= 64'h168b6f0d63a984c4;
        9'h12e: val <= 64'h257c729bc7b4c87e;
        9'h12f: val <= 64'h3f9503868ac974cb;
        9'h130: val <= 64'hcb6dff42caa0f1dd;
        9'h131: val <= 64'h31946bcd1b16766c;
        9'h132: val <= 64'h2e8539d6bafe5da0;
        9'h133: val <= 64'ha9fab3f584b6442f;
        9'h134: val <= 64'h304d13b1dc67994e;
        9'h135: val <= 64'he34623402e2f8494;
        9'h136: val <= 64'h2ee58b8ae5f3b86a;
        9'h137: val <= 64'he2a06c2b1ceacd85;
        9'h138: val <= 64'h406b21807c777ddd;
        9'h139: val <= 64'he3e3921cb82d869f;
        9'h13a: val <= 64'h5ce132b29b6d73d2;
        9'h13b: val <= 64'hb9b5f5173deee6cc;
        9'h13c: val <= 64'h28a75704b6f832a5;
        9'h13d: val <= 64'h8ab290a59fe3cfc0;
        9'h13e: val <= 64'hfc7ef36bab111162;
        9'h13f: val <= 64'h6967f31781645119;
        9'h140: val <= 64'ha45f1af7d2245cb9;
        9'h141: val <= 64'hbc3acebf6b9c2b5b;
        9'h142: val <= 64'h8e298479c0a0e66b;
        9'h143: val <= 64'h87b5dbaf841d059b;
        9'h144: val <= 64'h81bd00b0de2c9d82;
        9'h145: val <= 64'hc0d3b7deffa77d5a;
        9'h146: val <= 64'h02a3df308f452448;
        9'h147: val <= 64'h8b7b05e1ca3981c0;
        9'h148: val <= 64'hc417df5e89f7b642;
        9'h149: val <= 64'hb73d34f2df934901;
        9'h14a: val <= 64'h8663d3a47497698c;
        9'h14b: val <= 64'ha3a62eb9275e35bf;
        9'h14c: val <= 64'h167922d649cb9882;
        9'h14d: val <= 64'h7f351818f1790af8;
        9'h14e: val <= 64'h30f8aa43fbba9541;
        9'h14f: val <= 64'hb5ad86df652b9c54;
        9'h150: val <= 64'ha4e5d215de3b80da;
        9'h151: val <= 64'h9701ac7fd901b641;
        9'h152: val <= 64'hc1573945593890d3;
        9'h153: val <= 64'h4a92a0380919f7d1;
        9'h154: val <= 64'h7a36717da7661215;
        9'h155: val <= 64'h425d920eb06e0042;
        9'h156: val <= 64'hd381fa010bcc9a9f;
        9'h157: val <= 64'h713b005041fc3c82;
        9'h158: val <= 64'h04d3d5b73f71eeab;
        9'h159: val <= 64'h3574bf1c917a3610;
        9'h15a: val <= 64'h5bf09316ef57aba2;
        9'h15b: val <= 64'h4548bd13b03368aa;
        9'h15c: val <= 64'h04cf2c6d6cce4192;
        9'h15d: val <= 64'h6b57aa53e5a98d70;
        9'h15e: val <= 64'h1d9b90d76b42f0c9;
        9'h15f: val <= 64'h7da41c3873de1ff4;
        9'h160: val <= 64'h0387b4f2751bd978;
        9'h161: val <= 64'h175f0764d4fe699d;
        9'h162: val <= 64'hd527d7962f7f022b;
        9'h163: val <= 64'hd5db27b70d0b135c;
        9'h164: val <= 64'hbd3ec23314b2cd56;
        9'h165: val <= 64'h5efa891ff6dbaf67;
        9'h166: val <= 64'h3bcf449f234b5891;
        9'h167: val <= 64'hdbc63d905febe137;
        9'h168: val <= 64'h06116d6e36d122a8;
        9'h169: val <= 64'h920113e3af79396d;
        9'h16a: val <= 64'hc2f35829c95d6453;
        9'h16b: val <= 64'h93df7261d605955a;
        9'h16c: val <= 64'ha79726ec871e1065;
        9'h16d: val <= 64'hf47202a7a50bec5a;
        9'h16e: val <= 64'ha85c3659d43de854;
        9'h16f: val <= 64'h928536f96d4ea1c3;
        9'h170: val <= 64'h924a8af9f1b579a4;
        9'h171: val <= 64'h7a5a6636fff4d8d5;
        9'h172: val <= 64'hc40b456cc97a724a;
        9'h173: val <= 64'hecb1d5b1288c0467;
        9'h174: val <= 64'h2828695efb47245c;
        9'h175: val <= 64'h868c26d82900cb9f;
        9'h176: val <= 64'h320925fb60dbfe8e;
        9'h177: val <= 64'h54867c27853eea50;
        9'h178: val <= 64'h168afd615af96015;
        9'h179: val <= 64'hbdfe992cbe856aae;
        9'h17a: val <= 64'h7275817ef15ba564;
        9'h17b: val <= 64'hb8d5d7e2b0bb27cf;
        9'h17c: val <= 64'h0952740a0b6842ac;
        9'h17d: val <= 64'h46cf1fcf791e674b;
        9'h17e: val <= 64'ha62d5656acd524b6;
        9'h17f: val <= 64'hff2c61803344d752;
        9'h180: val <= 64'h7d88693cbcd06c09;
        9'h181: val <= 64'hc1c144299cfad4db;
        9'h182: val <= 64'hf285ae27eaa18986;
        9'h183: val <= 64'h2096da01cb0e1395;
        9'h184: val <= 64'h1411a00e391b2b05;
        9'h185: val <= 64'hf031a3c837e93bee;
        9'h186: val <= 64'h1613ab5002376e95;
        9'h187: val <= 64'h533fcc3337f034d6;
        9'h188: val <= 64'h699e09e27fb5a2f7;
        9'h189: val <= 64'hba7800393227d63e;
        9'h18a: val <= 64'heb396a20f99286dc;
        9'h18b: val <= 64'hbbd6285dbf40d56e;
        9'h18c: val <= 64'haa766d62016c2d11;
        9'h18d: val <= 64'h5b34bdac2ffe968b;
        9'h18e: val <= 64'hd30a7261a8061347;
        9'h18f: val <= 64'h917e98d79b317715;
        9'h190: val <= 64'h8bb73165987af370;
        9'h191: val <= 64'hd5c545c682869f5e;
        9'h192: val <= 64'h841f84c13becddb2;
        9'h193: val <= 64'hd4afb70e44bba9ae;
        9'h194: val <= 64'h8c108dbe401b459d;
        9'h195: val <= 64'h6076c43f94788282;
        9'h196: val <= 64'hb636cc24e8bf20f7;
        9'h197: val <= 64'hc224f984a0b324df;
        9'h198: val <= 64'h3e6f11b803888f52;
        9'h199: val <= 64'hc165e2c1105545d3;
        9'h19a: val <= 64'h7bb7ebfb3bd7e96e;
        9'h19b: val <= 64'h10e0d49b3864a97a;
        9'h19c: val <= 64'h52508c7d38d7ba63;
        9'h19d: val <= 64'hfdce873f04b3cdcf;
        9'h19e: val <= 64'ha774902ec6c71c46;
        9'h19f: val <= 64'hb67866d7b4a365e7;
        9'h1a0: val <= 64'hf7b4ba2d9df0d5c0;
        9'h1a1: val <= 64'he0635bd0b93a1bdc;
        9'h1a2: val <= 64'h0c4a7fbe051ff398;
        9'h1a3: val <= 64'hf87c8efe4b6288bf;
        9'h1a4: val <= 64'h78fc1fbb4bcf500a;
        9'h1a5: val <= 64'h4bdee7be591d901b;
        9'h1a6: val <= 64'h0b1e865068d7b92f;
        9'h1a7: val <= 64'h3c21dfe9964aa27d;
        9'h1a8: val <= 64'h69cc2499b5d0e006;
        9'h1a9: val <= 64'hd62c8b0f0163a483;
        9'h1aa: val <= 64'hecd30f2c264283c9;
        9'h1ab: val <= 64'h433e2054c542a8d9;
        9'h1ac: val <= 64'h7e2cf78941c21b7d;
        9'h1ad: val <= 64'h8b55fd4f7f43093e;
        9'h1ae: val <= 64'h2f8fe88b39eb0424;
        9'h1af: val <= 64'hfe520b7d0d189b15;
        9'h1b0: val <= 64'h945cad3144e4447b;
        9'h1b1: val <= 64'had96d27b765b2e07;
        9'h1b2: val <= 64'hac53caf7f8c7a080;
        9'h1b3: val <= 64'hd5f94fb789fcc0b5;
        9'h1b4: val <= 64'hf40c3c663d06f967;
        9'h1b5: val <= 64'h465a5076e16617d4;
        9'h1b6: val <= 64'h6eda213545239dda;
        9'h1b7: val <= 64'had04af2dd0a5cdf8;
        9'h1b8: val <= 64'h6c0a05cf5fcc99f4;
        9'h1b9: val <= 64'h5eb2e1219532b462;
        9'h1ba: val <= 64'h834dcee93a607d01;
        9'h1bb: val <= 64'h89f54d8aca46877e;
        9'h1bc: val <= 64'h281df540be5d6dc6;
        9'h1bd: val <= 64'h28edcd781a64dff0;
        9'h1be: val <= 64'hd9e7ea079a9837ae;
        9'h1bf: val <= 64'hc200c34c428c0ab7;
        9'h1c0: val <= 64'hebe7a64e376b5830;
        9'h1c1: val <= 64'h298f2a16e3a4ed08;
        9'h1c2: val <= 64'h0c53fe4b13b112c6;
        9'h1c3: val <= 64'haa67b391acc3ef09;
        9'h1c4: val <= 64'h18f502cda3c28201;
        9'h1c5: val <= 64'hd4290eefa37a465d;
        9'h1c6: val <= 64'h428c690577b9c856;
        9'h1c7: val <= 64'h2b21d5d29b29fc48;
        9'h1c8: val <= 64'hcab5591872b7e204;
        9'h1c9: val <= 64'hed4ef0482a20a18c;
        9'h1ca: val <= 64'hc00fc39c63e7f966;
        9'h1cb: val <= 64'h0e09bc1e8dde8e94;
        9'h1cc: val <= 64'h9d710fa0ed8c24ae;
        9'h1cd: val <= 64'h62d8f9ae5b30dc66;
        9'h1ce: val <= 64'h72f50c2cbafab647;
        9'h1cf: val <= 64'hbcbc6ef0d6fc3056;
        9'h1d0: val <= 64'h29de87ef8f67d937;
        9'h1d1: val <= 64'h38223fa950ae6665;
        9'h1d2: val <= 64'h0d22323b7caf731e;
        9'h1d3: val <= 64'h073186b31538a418;
        9'h1d4: val <= 64'hbaeac489f5800ccd;
        9'h1d5: val <= 64'h6cb3069e8edb6804;
        9'h1d6: val <= 64'hd76d203f8d07fd66;
        9'h1d7: val <= 64'h4f09b06851f19b8c;
        9'h1d8: val <= 64'h1da05a2f9a50479c;
        9'h1d9: val <= 64'ha3e301bf02afc0d3;
        9'h1da: val <= 64'hc16b84e71c229cc8;
        9'h1db: val <= 64'h5c2000d252a65e13;
        9'h1dc: val <= 64'hbad4e8a689f46332;
        9'h1dd: val <= 64'hac9b55f2101e876a;
        9'h1de: val <= 64'h65cf78db2da273fe;
        9'h1df: val <= 64'ha4585fce34d2787b;
        9'h1e0: val <= 64'h88ca46a8db06ac41;
        9'h1e1: val <= 64'h710ffc729d2eb8bb;
        9'h1e2: val <= 64'hb26d59578e5ff1f4;
        9'h1e3: val <= 64'h50fe397aab3b3c01;
        9'h1e4: val <= 64'h9d389e2168aa586c;
        9'h1e5: val <= 64'haab43810d00a3eef;
        9'h1e6: val <= 64'h4b3fa65af7dea24b;
        9'h1e7: val <= 64'h8242589591975ac5;
        9'h1e8: val <= 64'hd57f43ffda8d0c17;
        9'h1e9: val <= 64'h3983c4455e4f7165;
        9'h1ea: val <= 64'h3c3f1a77d7802a27;
        9'h1eb: val <= 64'h76b9f40e6a8cfd7a;
        9'h1ec: val <= 64'h60dbbd52adf1024d;
        9'h1ed: val <= 64'hfd7d962b2b5fac3d;
        9'h1ee: val <= 64'h2fcc31d52f27c41d;
        9'h1ef: val <= 64'h348243316172d144;
        9'h1f0: val <= 64'h51bbd36400249c33;
        9'h1f1: val <= 64'ha82ee1802e716e73;
        9'h1f2: val <= 64'h17f9860a7fdd34c6;
        9'h1f3: val <= 64'h9e636b690e69dfa4;
        9'h1f4: val <= 64'h97d0d4aadb3ca6ea;
        9'h1f5: val <= 64'h02701decf509064b;
        9'h1f6: val <= 64'h55c9ddc82171aeec;
        9'h1f7: val <= 64'ha1eeb77d1e63b2ef;
        9'h1f8: val <= 64'h6ec563543c68d9f8;
        9'h1f9: val <= 64'he19f42395d518aad;
        9'h1fa: val <= 64'h52a87a5cd4f7ad5e;
        9'h1fb: val <= 64'h07b3abdade355c36;
        9'h1fc: val <= 64'heebae03b172498fa;
        9'h1fd: val <= 64'hdc2abddc61622a91;
        9'h1fe: val <= 64'h84c0cccbc5ce6d1b;
        default: val <= 0;
    endcase
end

endmodule
